//--------------------------------------
//Project: The UVM environemnt for RegisterRTL
//Function: Register Config Transaction
//Author:  Le Hoang Van
//Page:    VLSI Technology
//--------------------------------------

// RegConfig Interface
interface RegConfig_Interface;
  // Content
endinterface: RegConfig_Interface
