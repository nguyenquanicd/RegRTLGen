//--------------------------------------
//Project: The UVM environemnt for RegisterRTL
//Function: Register Config Interface
//Author:  Nguyen Hung Quan, Le Hoang Van, Le Tan Thinh
//Page:    VLSI Technology
//--------------------------------------

interface RegConfig_Interface;
  // Content
endinterface: RegConfig_Interface
